module main

import credits

fn main() {
	credits.print_credits()
}
